
module modulo_uno (input INTERRUPTOR, output led );

    assign led = INTERRUPTOR;
endmodule